----------------------------------------------------------------------------------
-- Author: Stephan Proß
--
-- Create Date: 03/08/2022 02:46:11 PM
-- Design Name:
-- Module Name: Sorter Template
-- Project Name: BitSerialCompareSwap
-- Tool Versions: Vivado 2021.2
--
----------------------------------------------------------------------------------

library IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.NUMERIC_STD.all;

library work;
  use work.CustomTypes.all;

entity SORTER is
  generic (
    -- Bit-width of words
    W     : integer := 8;
    -- Number of input words.
    N     : integer := 4;
    -- Number of sorted ouput words.
    M     : integer := 4;
    -- Number of available BRAMs
    NUM_BRAM : integer := 4

  );
  port (
    -- System clock
    CLK          : in    std_logic;
    -- Enable signal
    E            : in    std_logic;
    -- Syncronous reset
    RST          : in    std_logic;
    -- Parallel input of N unsorted w-bit words.
    PAR_INPUT    : in    SLVArray(0 to N - 1)(W-1 downto 0);
    -- Parallel ouput of N sorted w-bit words.
    PAR_OUTPUT   : out   SLVArray(0 to M - 1)(W-1 downto 0)
  );
end entity SORTER;

architecture STRUCTURAL of SORTER is
  -- Number of BRAM blocks required per IO.
  constant BRAM_PER_IO : integer := (W + 32 - 1) / 32;
  -- Number of available IO ports replacable with BRAM version.
  constant NUM_IO_BRAM : integer := NUM_BRAM / BRAM_PER_IO;

  -- Number of remaining BRAMS for output deserialization.
  constant NUM_OUTPUT_BRAM : integer := NUM_IO_BRAM - N;

  -- Start signal generated by cycle timer.
  signal start_i      : std_logic;
  -- Done signal generated by the sorting network.
  signal done_i       : std_logic;
  -- Serial unsorted data.
  signal ser_unsorted_i  : std_logic_vector(0 to N - 1);
  -- Serial sorted data.
  signal ser_sorted_i : std_logic_vector(0 to M - 1);

begin

  CYCLE_TIMER_1 : entity work.cycle_timer
    generic map (
      W => W,
      DELAY => 0
    )
    port map (
      CLK   => CLK,
      RST   => RST,
      E     => E,
      START => start_i
    );

  IO_SERIZALIZERS_MIXED : if (N > NUM_IO_BRAM) generate

    -- Fill the remainder of required serializers with shift-register variants.
    SERIALIZER_BRAM_1 : entity work.serializer_bram
      generic map (
        N => NUM_IO_BRAM ,
        W => W
      )
      port map (
        CLK        => CLK,
        RST        => RST,
        E          => E,
        LOAD       => start_i,
        PAR_INPUT  => PAR_INPUT(0 to NUM_IO_BRAM-1),
        SER_OUTPUT => ser_unsorted_i(0 to NUM_IO_BRAM-1)
      );

    SERIALIZER_SR_1 : entity work.serializer_sr
      generic map (
        N => N - NUM_IO_BRAM ,
        W => W
      )
      port map (
        CLK        => CLK,
        RST        => RST,
        E          => E,
        LOAD       => start_i,
        PAR_INPUT  => PAR_INPUT(NUM_IO_BRAM to N-1),
        SER_OUTPUT => ser_unsorted_i(NUM_IO_BRAM to N -1)
      );

  end generate IO_SERIZALIZERS_MIXED;

  IO_SERIALIZERS_BRAM : if (N <= NUM_IO_BRAM) generate

    -- We can use only BRAM serializers for input.
    SERIALIZER_BRAM_2 : entity work.serializer_bram
      generic map (
        N => N,
        W => W
      )
      port map (
        CLK        => CLK,
        RST        => RST,
        E          => E,
        LOAD       => start_i,
        PAR_INPUT  => PAR_INPUT,
        SER_OUTPUT => ser_unsorted_i
      );

 end generate IO_SERIALIZERS_BRAM;

  IO_SERIALIZERS_SR : if (NUM_IO_BRAM = 0) generate

    -- There is no BRAM available for serialization.
    SERIALIZER_SR_2 : entity work.serializer_SR
      generic map (
        N => N,
        W => W
      )
      port map (
        CLK        => CLK,
        RST        => RST,
        E          => E,
        LOAD       => start_i,
        PAR_INPUT  => PAR_INPUT,
        SER_OUTPUT => ser_unsorted_i
      );

 end generate IO_SERIALIZERS_SR;

  SORTING_NETWORK_1 : entity work.oddeven_4_to_4_max
    generic map (
      W => W
    )
    port map (
      CLK        => CLK,
      RST        => RST,
      E          => E,
      START      => start_i,
      SER_INPUT  => ser_unsorted_i,
      DONE       => done_i,
      SER_OUTPUT => ser_sorted_i
    );

  IO_DESERIZALIZERS_MIXED : if (M > NUM_OUTPUT_BRAM and NUM_OUTPUT_BRAM > 0) generate

    -- Fill the remainder of required deserializers with shift-register variants.
    DESERIALIZER_BRAM_1 : entity work.deserializer_bram
      generic map (
        N => NUM_OUTPUT_BRAM,
        W => W
      )
      port map (
        CLK        => CLK,
        RST        => RST,
        E          => E,
        STORE      => done_i,
        SER_INPUT  => ser_sorted_i(0 to NUM_OUTPUT_BRAM-1),
        PAR_OUTPUT => PAR_OUTPUT(0 to NUM_OUTPUT_BRAM -1)
      );

    DESERIALIZER_SR_1 : entity work.deserializer_sr
      generic map (
        N => M - NUM_OUTPUT_BRAM,
        W => W
      )
      port map (
        CLK        => CLK,
        RST        => RST,
        E          => E,
        STORE      => done_i,
        SER_INPUT  => ser_sorted_i(NUM_OUTPUT_BRAM to M - 1),
        PAR_OUTPUT => PAR_OUTPUT(NUM_OUTPUT_BRAM to M - 1)
      );

    end generate IO_DESERIZALIZERS_MIXED;

  IO_DESERIZALIZERS_BRAM : if (M <= NUM_OUTPUT_BRAM and NUM_OUTPUT_BRAM > 0) generate

    -- We have enough BRAMs for the entire output.
    DESERIALIZER_BRAM_2 : entity work.deserializer_bram
      generic map (
        N => M,
        W => W
      )
      port map (
        CLK        => CLK,
        RST        => RST,
        E          => E,
        STORE      => done_i,
        SER_INPUT  => ser_sorted_i,
        PAR_OUTPUT => PAR_OUTPUT
      );

  end generate IO_DESERIZALIZERS_BRAM;

  IO_DESERIZALIZERS_SR : if (NUM_OUTPUT_BRAM <= 0) generate

    -- There are no available BRAMs for output deserialization.
    DESERIALIZER_SR_2 : entity work.deserializer_sr
      generic map (
        N => M,
        W => W
      )
      port map (
        CLK        => CLK,
        RST        => RST,
        E          => E,
        STORE      => done_i,
        SER_INPUT  => ser_sorted_i,
        PAR_OUTPUT => PAR_OUTPUT
      );

  end generate IO_DESERIZALIZERS_SR;
end architecture STRUCTURAL;
